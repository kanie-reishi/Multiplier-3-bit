library verilog;
use verilog.vl_types.all;
entity mul3Bit_vlg_vec_tst is
end mul3Bit_vlg_vec_tst;
