library verilog;
use verilog.vl_types.all;
entity mul3Bit_vlg_check_tst is
    port(
        S               : in     vl_logic_vector(5 downto 0);
        sampler_rx      : in     vl_logic
    );
end mul3Bit_vlg_check_tst;
